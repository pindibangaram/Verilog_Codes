module up_down_8bit_tb();
  reg clk,rst,load,updown;
  reg [7:0]data_in;
  wire [7:0]count;
  
